../chisel/verilog/ofdm_demodulator.v